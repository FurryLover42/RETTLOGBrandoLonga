library ieee;
use ieee.std_logic_1164.all;

--	The syntax for an entity with a port in VHDL is:
--	entity <entity_name> is
--	port(
--	    <entity_signal_name> : in|out|inout <signal_type>;
--	    ...
--	);
--	end entity;
--	
--	The syntax for instantiating such a module in another VHDL file is:
--	<label> : entity <library_name>.<entity_name>(<architecture_name>) port map(
--	    <entity_signal_name> => <local_signal_name>,
--	    ...
--	);
--	
--	The <label> can be any name, and it will show up in the hierarchy window in ModelSim.
--	The <library_name> for a module is set in the simulator, not in the VHDL code. By default every module is compiled into the work library.
--	The <entity_name> and <architecture_name> must match the module we are creating an instance of.
--	Finally, each of the entity signals must be mapped to a local signal name.




entity fsm_tb is	
end fsm_tb;


architecture sim of fsm_tb is

	signal input:	std_logic;
	signal clk:		std_logic;
	signal reset:	std_logic;
	signal output:	std_logic;

begin
	
	--port mapping
	finite_state_machine : entity work.fsm(rtl) port map(
		input	=> input,
		clk		=> clk,
		reset	=> reset,
		output	=> output);
	
	--clock process
	process is
	begin
		clk <= '0';
		wait for 10 ns;
		clk <= '1';
		wait for 10 ns;
	end process;
	
	--testbench process
	process is
	begin
		input <= '0';
		reset <= '1';
		wait for 28 ns;
		reset <= '0';
		input <= '1';
		wait for 85 ns;
		input <= '0';
		wait for 20 ns;
		input <= '1';
		wait for 23 ns;
		input <= '0';
		wait for 30 ns;
		input <= '1';
		wait for 7 ns;
		input <= '0';
		wait for 23 ns;
		input <= '1';
		wait for 12 ns;
		input <= '0';
		wait for 19 ns;
		input <= '1';
		wait for 10 ns;
		input <= '0';
		wait for 13 ns;
		input <= '1';
		wait for 29 ns;
		input <= '0';
		wait for 10 ns;
		input <= '1';
		wait for 90 ns;
		input <= '0';
		wait for 20 ns;
		input <= '1';
		wait for 94 ns;
		reset <= '1';
		wait for 55 ns;
		input <= '0';
		reset <= '0';
		wait for 24 ns;
		input <= '1';
		wait;
		
	end process;
	

end architecture sim;
-- va bene anche solo end sim;